module pc_vga_8x16_80_FF (
	 input		clk,
	 input  [6:0]	ascii_code,
	 input  [3:0]	row,
	 input  [2:0]  col,
	 output wire	row_of_pixels
	 );

RAMB16_S1 BRAM_PC_VGA_0 (
	.CLK(clk),
	.EN(1'b1),
	.WE(1'b0),
	.ADDR({ascii_code[6:1], ~ascii_code[0], row, ~col}),
	.SSR(1'b0),
	.DI(1'b0),
	.DO(row_of_pixels)
	);
	 
defparam BRAM_PC_VGA_0.INIT_00 = 256'h00007c060c3c66c2c0c0c0c2663c00000000000076cccccccccccc0000cc0000;
defparam BRAM_PC_VGA_0.INIT_01 = 256'h000000007cc6c0c0fec67c0030180c000000000076cccccc7c0c78006c381000;
defparam BRAM_PC_VGA_0.INIT_02 = 256'h0000000076cccccc7c0c780000cc00000000000076cccccc7c0c780018306000;
defparam BRAM_PC_VGA_0.INIT_03 = 256'h0000000076cccccc7c0c7800386c38000000003c060c3c666060663c00000000;
defparam BRAM_PC_VGA_0.INIT_04 = 256'h000000007cc6c0c0fec67c006c381000000000007cc6c0c0fec67c0000c60000;
defparam BRAM_PC_VGA_0.INIT_05 = 256'h000000007cc6c0c0fec67c0018306000000000003c1818181818380000660000;
defparam BRAM_PC_VGA_0.INIT_06 = 256'h000000003c18181818183800663c1800000000003c1818181818380018306000;
defparam BRAM_PC_VGA_0.INIT_07 = 256'h00000000c6c6c6fec6c66c381000c60000000000c6c6c6fec6c66c3800386c38;
defparam BRAM_PC_VGA_0.INIT_08 = 256'h00000000fe6660607c6066fe006030180000000077dcd87e1b3b6e0000000000;
defparam BRAM_PC_VGA_0.INIT_09 = 256'h00000000ceccccccccfecccc6c3e0000000000007cc6c6c6c6c67c006c381000;
defparam BRAM_PC_VGA_0.INIT_0A = 256'h000000007cc6c6c6c6c67c0000c60000000000007cc6c6c6c6c67c0018306000;
defparam BRAM_PC_VGA_0.INIT_0B = 256'h0000000076cccccccccccc00cc7830000000000076cccccccccccc0018306000;
defparam BRAM_PC_VGA_0.INIT_0C = 256'h00780c067ec6c6c6c6c6c60000c60000000000007cc6c6c6c6c6c6c67c00c600;
defparam BRAM_PC_VGA_0.INIT_0D = 256'h000000007cc6c6c6c6c6c6c6c600c6000000000018187ec3c0c0c0c37e181800;
defparam BRAM_PC_VGA_0.INIT_0E = 256'h00000000fce660606060f060646c380000000000181818ff18ff183c66c30000;
defparam BRAM_PC_VGA_0.INIT_0F = 256'h00000000f36666666f66627c6666fc00000070d818181818187e1818181b0e00;

defparam BRAM_PC_VGA_0.INIT_10 = 256'h0000000076cccccc7c0c780060301800000000003c1818181818380030180c00;
defparam BRAM_PC_VGA_0.INIT_11 = 256'h000000007cc6c6c6c6c67c00603018000000000076cccccccccccc0060301800;
defparam BRAM_PC_VGA_0.INIT_12 = 256'h00000000666666666666dc00dc76000000000000c6c6c6cedefef6e6c600dc76;
defparam BRAM_PC_VGA_0.INIT_13 = 256'h0000000000000000007e003e6c6c3c000000000000000000007c00386c6c3800;
defparam BRAM_PC_VGA_0.INIT_14 = 256'h000000007cc6c6c060303000303000000000000000c0c0c0c0fe000000000000;
defparam BRAM_PC_VGA_0.INIT_15 = 256'h000000000006060606fe00000000000000001f0c069bce603018ccc6c2c0c000;
defparam BRAM_PC_VGA_0.INIT_16 = 256'h000006063e96ce663018ccc6c2c0c00000000000183c3c3c1818180018180000;
defparam BRAM_PC_VGA_0.INIT_17 = 256'h000000000000366cd86c360000000000000000000000d86c366cd80000000000;
defparam BRAM_PC_VGA_0.INIT_18 = 256'h44114411441144114411441144114411aa55aa55aa55aa55aa55aa55aa55aa55;
defparam BRAM_PC_VGA_0.INIT_19 = 256'h77dd77dd77dd77dd77dd77dd77dd77dd18181818181818181818181818181818;
defparam BRAM_PC_VGA_0.INIT_1A = 256'h1818181818181818f8181818181818181818181818181818f818f81818181818;
defparam BRAM_PC_VGA_0.INIT_1B = 256'h3636363636363636f6363636363636363636363636363636fe00000000000000;
defparam BRAM_PC_VGA_0.INIT_1C = 256'h1818181818181818f818f800000000003636363636363636f606f63636363636;
defparam BRAM_PC_VGA_0.INIT_1D = 256'h363636363636363636363636363636363636363636363636f606fe0000000000;
defparam BRAM_PC_VGA_0.INIT_1E = 256'h0000000000000000fe06f636363636360000000000000000fe36363636363636;
defparam BRAM_PC_VGA_0.INIT_1F = 256'h0000000000000000f818f818181818181818181818181818f800000000000000;

defparam BRAM_PC_VGA_0.INIT_20 = 256'h00000000000000001f181818181818180000000000000000ff18181818181818;
defparam BRAM_PC_VGA_0.INIT_21 = 256'h1818181818181818ff0000000000000018181818181818181f18181818181818;
defparam BRAM_PC_VGA_0.INIT_22 = 256'h0000000000000000ff000000000000001818181818181818ff18181818181818;
defparam BRAM_PC_VGA_0.INIT_23 = 256'h18181818181818181f181f181818181836363636363636363736363636363636;
defparam BRAM_PC_VGA_0.INIT_24 = 256'h00000000000000003f30373636363636363636363636363637303f0000000000;
defparam BRAM_PC_VGA_0.INIT_25 = 256'h0000000000000000ff00f736363636363636363636363636f700ff0000000000;
defparam BRAM_PC_VGA_0.INIT_26 = 256'h363636363636363637303736363636360000000000000000ff00ff0000000000;
defparam BRAM_PC_VGA_0.INIT_27 = 256'h3636363636363636f700f736363636360000000000000000ff00ff1818181818;
defparam BRAM_PC_VGA_0.INIT_28 = 256'h0000000000000000ff363636363636361818181818181818ff00ff0000000000;
defparam BRAM_PC_VGA_0.INIT_29 = 256'h3636363636363636ff0000000000000000000000000000003f36363636363636;
defparam BRAM_PC_VGA_0.INIT_2A = 256'h00000000000000001f181f181818181818181818181818181f181f0000000000;
defparam BRAM_PC_VGA_0.INIT_2B = 256'h36363636363636363f000000000000003636363636363636ff36363636363636;
defparam BRAM_PC_VGA_0.INIT_2C = 256'h1818181818181818ff18ff18181818180000000000000000f818181818181818;
defparam BRAM_PC_VGA_0.INIT_2D = 256'h18181818181818181f00000000000000ffffffffffffffffffffffffffffffff;
defparam BRAM_PC_VGA_0.INIT_2E = 256'hffffffffffffffffff00000000000000f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0;
defparam BRAM_PC_VGA_0.INIT_2F = 256'h0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f000000000000000000ffffffffffffff;

defparam BRAM_PC_VGA_0.INIT_30 = 256'h0000000076dcd8d8d8dc76000000000000000000ccc6c6c6ccd8cccccc780000;
defparam BRAM_PC_VGA_0.INIT_31 = 256'h00000000c0c0c0c0c0c0c0c6c6fe0000000000006c6c6c6c6c6c6cfe00000000;
defparam BRAM_PC_VGA_0.INIT_32 = 256'h00000000fec66030183060c6fe0000000000000070d8d8d8d8d87e0000000000;
defparam BRAM_PC_VGA_0.INIT_33 = 256'h000000c060607c66666666660000000000000000181818181818dc7600000000;
defparam BRAM_PC_VGA_0.INIT_34 = 256'h000000007e183c6666663c187e00000000000000386cc6c6fec6c66c38000000;
defparam BRAM_PC_VGA_0.INIT_35 = 256'h00000000ee6c6c6c6cc6c6c66c380000000000003c666666663e0c18301e0000;
defparam BRAM_PC_VGA_0.INIT_36 = 256'h0000000000007edbdbdb7e000000000000000000c0607ef3dbdb7e0603000000;
defparam BRAM_PC_VGA_0.INIT_37 = 256'h000000001c306060607c6060301c000000000000c6c6c6c6c6c6c6c67c000000;
defparam BRAM_PC_VGA_0.INIT_38 = 256'h0000000000fe0000fe0000fe0000000000000000ff000018187e181800000000;
defparam BRAM_PC_VGA_0.INIT_39 = 256'h000000007e0030180c060c1830000000000000007e000c18306030180c000000;
defparam BRAM_PC_VGA_0.INIT_3A = 256'h181818181818181818181b1b1b0e00000000000070d8d8d81818181818181818;
defparam BRAM_PC_VGA_0.INIT_3B = 256'h00000000001818007e00181800000000000000000000dc7600dc760000000000;
defparam BRAM_PC_VGA_0.INIT_3C = 256'h0000000000000000000000386c6c380000000000000000181800000000000000;
defparam BRAM_PC_VGA_0.INIT_3D = 256'h00000000000000180000000000000000000000001c3c6c6cec0c0c0c0c0c0f00;
defparam BRAM_PC_VGA_0.INIT_3E = 256'h0000000000000000006c6c6c6c6cd800000000000000000000f8c86030d87000;
defparam BRAM_PC_VGA_0.INIT_3F = 256'h00000000007c7c7c7c7c7c7c0000000000000000000000000000000000000000;
	 
endmodule
